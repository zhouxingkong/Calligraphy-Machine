/*
��ģ��Ĺ�������֤ʵ�ֺ�PC�����л����Ĵ���ͨ�ŵĹ��ܡ���Ҫ��PC���ϰ�װһ�����ڵ��Թ�������֤����Ĺ��ܡ�
����ʵ����һ���շ�һ֡10��bit��������żУ��λ���Ĵ��ڿ�������10��bit��1λ��ʼλ��8������λ��1������λ��
���ڵĲ������ɳ����ж����div_par�������������ĸò�������ʵ����Ӧ�Ĳ����ʡ�����ǰ�趨��div_par ��ֵ
��0x104����Ӧ�Ĳ�������9600����һ��8�������ʵ�ʱ�ӽ����ͻ����ÿһλbit������ʱ�仮��Ϊ8��ʱ϶��ʹͨ
��ͬ��.

����Ļ������������ǣ�����һ������SW0����������PC�Ĵ��ڷ��͡�welcome"��
PC�����պ���ʾ��֤�����Ƿ���ȷ�����ڵ��Թ�����ɰ�ASCII����ܷ�ʽ��.
PC����ʱ��CPLD����0-F��ʮ���������ݣ�CPLD���ܺ���ʾ��7���������.
*/
module serial(clk,rxd,txd,rxd_buf,rxd_ok,on
);

input clk;
input rxd;//�������ݽ���
output txd;//�������ݷ��Ͷ�
output reg[7:0] rxd_buf;//�������ݻ���
output reg rxd_ok=0;
input on;

//assign rxd_ok=(state_rec==4'd9||(state_rec==4'd0&&accept==0))?1:0;
wire rst=1;
////////////////////inner reg////////////////////
reg[15:0] div_reg;//��Ƶ����������Ƶֵ�ɲ����ʾ�������Ƶ��õ�Ƶ��8�������ʵ�ʱ��
reg[2:0]  div8_tras_reg;//�üĴ����ļ���ֵ��Ӧ����ʱ��ǰλ�ڵ�ʱ϶��
reg[2:0]  div8_rec_reg;//�üĴ����ļ���ֵ��Ӧ����ʱ��ǰλ�ڵ�ʱ϶��
reg[3:0] state_tras;//����״̬�Ĵ���
reg[3:0] state_rec;//����״̬�Ĵ���
reg clkbaud_tras;//�Բ�����ΪƵ�ʵķ���ʹ���ź�
reg clkbaud_rec;//�Բ�����ΪƵ�ʵĽ���ʹ���ź�
reg clkbaud8x;//��8��������ΪƵ�ʵ�ʱ�ӣ����������ǽ����ͻ����һ��bit��ʱ�����ڷ�Ϊ8��ʱ϶

reg recstart;//��ʼ���ͱ�־
reg recstart_tmp;

reg trasstart;//��ʼ���ܱ�־

reg rxd_reg1;//���ռĴ���1
reg rxd_reg2;//���ռĴ���2����Ϊ��������Ϊ�첽�źţ�������������
reg txd_reg;//���ͼĴ���

reg[7:0] txd_buf;//�������ݻ���

reg[2:0] send_state;//ÿ�ΰ�����PC����"Welcome"�ַ��������Ƿ���״̬�Ĵ���
reg[19:0] cnt_delay;//��ʱȥ��������
reg start_delaycnt;//��ʼ��ʱ������־
reg key_entry1,key_entry2;//ȷ���м����±�־

////////////////////////////////////////////////
parameter div_par=16'd651;//��Ƶ��������ֵ�ɶ�Ӧ�Ĳ����ʼ�����ã����˲�����Ƶ��ʱ��Ƶ���ǲ������ʵ�8	
		  //�����˴�ֵ��Ӧ9600�Ĳ����ʣ�����Ƶ����ʱ��Ƶ����9600*8

////////////////////////////////////////////////
assign txd=txd_reg;

always@(posedge clk )
begin
	if(!rst) begin 
		cnt_delay<=0;
		start_delaycnt<=0;
	 end
	else if(start_delaycnt) begin
		if(cnt_delay!=20'd800000) begin
			cnt_delay<=cnt_delay+1;
		 end
		else begin
			cnt_delay<=0;
			start_delaycnt<=0;
		 end
	 end
	else begin
		if(cnt_delay==0)
				start_delaycnt<=1;
	 end
end

always@(posedge clk)
begin
	if(!rst) 
		key_entry1<=0;
	else begin
		if(key_entry2)
			key_entry1<=0;
		else if(cnt_delay==20'd800000) begin
				key_entry1<=1;
		 end
	 end
end

always@(posedge clk )
begin
	if(!rst)
		div_reg<=0;
	else begin
		if(div_reg==div_par-1)
			div_reg<=0;
		else
			div_reg<=div_reg+1;
	 end
end

always@(posedge clk)//��Ƶ�õ�8�������ʵ�ʱ��
begin
	if(!rst)
		clkbaud8x<=0;
	else if(div_reg==div_par-1)
		clkbaud8x<=~clkbaud8x;
end


always@(posedge clkbaud8x or negedge rst)
begin
	if(!rst)
		div8_rec_reg<=0;
	else if(recstart)//���տ�ʼ��־
		div8_rec_reg<=div8_rec_reg+1;//���տ�ʼ��ʱ϶����8�������ʵ�ʱ���¼�1ѭ��
end

always@(posedge clkbaud8x or negedge rst)
begin
	if(!rst)
		div8_tras_reg<=0;
	else if(trasstart)
		div8_tras_reg<=div8_tras_reg+1;//���Ϳ�ʼ��ʱ϶����8�������ʵ�ʱ���¼�1ѭ��
end

always@(div8_rec_reg)
begin
	if(div8_rec_reg==7)
		clkbaud_rec=1;//�ڵ�7��ʱ϶������ʹ���ź���Ч�������ݴ���
	else
		clkbaud_rec=0;
end

always@(div8_tras_reg)
begin
	if(div8_tras_reg==7)
		clkbaud_tras=1;//�ڵ�7��ʱ϶������ʹ���ź���Ч�������ݷ���
	else
		clkbaud_tras=0;
end

always@(posedge clkbaud8x or negedge rst)
begin
	if(!rst) begin
		txd_reg<=1;
		trasstart<=0;
		txd_buf<=0;
		state_tras<=0;
		send_state<=0;
		key_entry2<=0;
	 end
	else begin
		if(!key_entry2) begin
			if(key_entry1) begin
				key_entry2<=1;
				txd_buf<=8'd119; //"w"
			 end
		 end
		else  begin
			case(state_tras)
				4'b0000: begin  //������ʼλ
					if(!trasstart&&send_state<7) 
						trasstart<=1;
					else if(send_state<7) begin
						if(clkbaud_tras) begin
							txd_reg<=0;
							state_tras<=state_tras+1;
						 end
					 end
					else begin
						key_entry2<=0;
						state_tras<=0;
					 end					
				end		
				4'b0001: begin //���͵�1λ
					if(clkbaud_tras) begin
						txd_reg<=txd_buf[0];
						txd_buf[6:0]<=txd_buf[7:1];
						state_tras<=state_tras+1;
					 end
				 end
				4'b0010: begin //���͵�2λ
					if(clkbaud_tras) begin
						txd_reg<=txd_buf[0];
						txd_buf[6:0]<=txd_buf[7:1];
						state_tras<=state_tras+1;
					 end
				 end
				 4'b0011: begin //���͵�3λ
				 	if(clkbaud_tras) begin
						txd_reg<=txd_buf[0];
						txd_buf[6:0]<=txd_buf[7:1];
						state_tras<=state_tras+1;
					 end
				 end
				4'b0100: begin //���͵�4λ
					if(clkbaud_tras) begin
						txd_reg<=txd_buf[0];
						txd_buf[6:0]<=txd_buf[7:1];
						state_tras<=state_tras+1;
					 end
				 end
				4'b0101: begin //���͵�5λ
					if(clkbaud_tras) begin
						txd_reg<=txd_buf[0];
						txd_buf[6:0]<=txd_buf[7:1];
						state_tras<=state_tras+1;
					 end
				 end
				4'b0110: begin //���͵�6λ
					if(clkbaud_tras) begin
						txd_reg<=txd_buf[0];
						txd_buf[6:0]<=txd_buf[7:1];
						state_tras<=state_tras+1;
					 end
				 end
				4'b0111: begin //���͵�7λ
					if(clkbaud_tras) begin
						txd_reg<=txd_buf[0];
						txd_buf[6:0]<=txd_buf[7:1];
						state_tras<=state_tras+1;
					 end
				 end
				4'b1000: begin //���͵�8λ
					if(clkbaud_tras) begin
						txd_reg<=txd_buf[0];
						txd_buf[6:0]<=txd_buf[7:1];
						state_tras<=state_tras+1;
					 end
				 end
				4'b1001: begin //����ֹͣλ
					if(clkbaud_tras) begin
						txd_reg<=1;
						txd_buf<=8'h55;
						state_tras<=state_tras+1;
					 end
				 end
				4'b1111:begin 
					if(clkbaud_tras) begin
						state_tras<=state_tras+1;
						send_state<=send_state+1;
						trasstart<=0;
						case(send_state)
							3'b000:
								txd_buf<=8'd101;//"e"
							3'b001:
								txd_buf<=8'd108;//"l"
							3'b010:
								txd_buf<=8'd99;//"c"
							3'b011:
								txd_buf<=8'd111;//"o"
							3'b100:
								txd_buf<=8'd109;//"m"
							3'b101:
								txd_buf<=8'd101;//"e"
							default:
								txd_buf<=0;
						 endcase
					 end
				 end
				default: begin
					if(clkbaud_tras) begin
						state_tras<=state_tras+1;
						trasstart<=1;
					 end
				 end
			 endcase
		 end
	 end
end

always@(posedge clkbaud8x or negedge rst)//����PC��������
begin
	if(!rst) begin
		rxd_reg1<=0;
		rxd_reg2<=0;
		rxd_buf<=0;
		state_rec<=0;
		recstart<=0;
		recstart_tmp<=0;
	 end
	else  begin
		 rxd_reg1<=rxd;
		 rxd_reg2<=rxd_reg1;
		 if(state_rec==0) begin
		      rxd_ok<=0;
			 if(recstart_tmp==1) begin
		 		recstart<=1;
		 		recstart_tmp<=0;
				state_rec<=state_rec+1;
		  	  end
		 	 else if(!rxd_reg1&&rxd_reg2) //��⵽��ʼλ���½��أ��������״̬
		 	    begin
				    recstart_tmp<=1;
				end
		   end
		 else if(state_rec>=1&&state_rec<=8) begin
		      rxd_ok<=0;
		 	 if(clkbaud_rec) begin
			 	rxd_buf[7]<=rxd_reg2;
				rxd_buf[6:0]<=rxd_buf[7:1];
				state_rec<=state_rec+1;
			  end
		  end
		 else if(state_rec==9) begin
		     rxd_ok<=1;
		 	 if(clkbaud_rec) begin
		 		state_rec<=10;
				recstart<=0;
			 end
		  end
		  else if(state_rec==10)begin
		      if(on==1) state_rec<=0;
		      else state_rec<=10;
		  end
	  end
end

endmodule
	
